module tb_fourBitSubtractor;
	reg [3:0] X, Y;
	wire [3:0] D;
	wire B;
	
	fourBitSubtractor UUT(X, Y, D, B);
	
	initial
		begin
			$dumpfile("tb_fourBitSubtractor.vpd");
			$dumpvars;
			
			// X = 4'd0; Y = 4'd0;
			// #10
			// X = 4'd1; Y = 4'd1;
			// #10
			// X = 4'd2; Y = 4'd2;
			// #10
			// X = 4'd3; Y = 4'd3;
			// #10
			// X = 4'd4; Y = 4'd4;
			// #10
			// X = 4'd5; Y = 4'd5;
			// #10
			// X = 4'd6; Y = 4'd6;
			// #10
			// X = 4'd7; Y = 4'd7;
			// #10
			// X = 4'd8; Y = 4'd8;
			// #10
			// X = 4'd9; Y = 4'd9;
			// #10
			// X = 4'd10; Y = 4'd10;
			// #10
			// X = 4'd11; Y = 4'd11;
			// #10
			// X = 4'd12; Y = 4'd12;
			// #10
			// X = 4'd13; Y = 4'd13;
			// #10
			// X = 4'd14; Y = 4'd14;
			// #10
			// X = 4'd15; Y = 4'd15;
			// #10
			
			X[3] = 1; X[2] = 0; X[1] = 1; X[0] = 0;
			Y[3] = 0; Y[2] = 1; Y[1] = 0; Y[0] = 1;
			#10
			
			X[3] = 1; X[2] = 1; X[1] = 0; X[0] = 1;
			Y[3] = 1; Y[2] = 0; Y[1] = 0; Y[0] = 0;
			#10
			
			X[3] = 0; X[2] = 1; X[1] = 0; X[0] = 0;
			Y[3] = 1; Y[2] = 1; Y[1] = 0; Y[0] = 0;
			#10
			
			X[3] = 1; X[2] = 1; X[1] = 1; X[0] = 1;
			Y[3] = 1; Y[2] = 1; Y[1] = 1; Y[0] = 0;
			#10
			
			X[3] = 0; X[2] = 0; X[1] = 1; X[0] = 0;
			Y[3] = 1; Y[2] = 0; Y[1] = 1; Y[0] = 0;
			#10
			
			X[3] = 1; X[2] = 1; X[1] = 1; X[0] = 1;
			Y[3] = 0; Y[2] = 1; Y[1] = 1; Y[0] = 1;
			#10
			
			X[3] = 0; X[2] = 1; X[1] = 1; X[0] = 0;
			Y[3] = 1; Y[2] = 0; Y[1] = 1; Y[0] = 0;
			#10
			
			X[3] = 1; X[2] = 1; X[1] = 0; X[0] = 1;
			Y[3] = 1; Y[2] = 1; Y[1] = 0; Y[0] = 1;
			#10
			
			X[3] = 1; X[2] = 0; X[1] = 0; X[0] = 0;
			Y[3] = 0; Y[2] = 1; Y[1] = 1; Y[0] = 0;
			#10
			
			X[3] = 1; X[2] = 0; X[1] = 1; X[0] = 0;
			Y[3] = 1; Y[2] = 1; Y[1] = 1; Y[0] = 1;
			#10
			
		$finish;
	end
endmodule