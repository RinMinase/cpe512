module tb_fourBitAdder;
	reg [3:0] X, Y;
	reg	Z;
	wire [3:0] S;
	wire C;
	
	fourBitAdder UUT(X, Y, Z, S, C);
	
	initial
		begin
			$dumpfile("tb_fourBitAdder.vpd");
			$dumpvars;
			
			// X = 4'd0; Y = 4'd0; Z = 0;
			// #10
			// X = 4'd1; Y = 4'd1; Z = 1;
			// #10
			// X = 4'd2; Y = 4'd2; Z = 0;
			// #10
			// X = 4'd3; Y = 4'd3; Z = 1;
			// #10
			// X = 4'd4; Y = 4'd4; Z = 0;
			// #10
			// X = 4'd5; Y = 4'd5; Z = 1;
			// #10
			// X = 4'd6; Y = 4'd6; Z = 0;
			// #10
			// X = 4'd7; Y = 4'd7; Z = 1;
			// #10
			// X = 4'd8; Y = 4'd8; Z = 0;
			// #10
			// X = 4'd9; Y = 4'd9; Z = 1;
			// #10
			// X = 4'd10; Y = 4'd10; Z = 0;
			// #10
			// X = 4'd11; Y = 4'd11; Z = 1;
			// #10
			// X = 4'd12; Y = 4'd12; Z = 0;
			// #10
			// X = 4'd13; Y = 4'd13; Z = 1;
			// #10
			// X = 4'd14; Y = 4'd14; Z = 0;
			// #10
			// X = 4'd15; Y = 4'd15; Z = 1;
			// #10

			X[3] = 1; X[2] = 0; X[1] = 1; X[0] = 0;
			Y[3] = 0; Y[2] = 1; Y[1] = 0; Y[0] = 1;
			Z = 0;
			#10
			
			X[3] = 1; X[2] = 1; X[1] = 0; X[0] = 1;
			Y[3] = 1; Y[2] = 0; Y[1] = 0; Y[0] = 0;
			Z = 1;
			#10
			
			X[3] = 0; X[2] = 1; X[1] = 0; X[0] = 0;
			Y[3] = 1; Y[2] = 1; Y[1] = 0; Y[0] = 0;
			Z = 0;
			#10
			
			X[3] = 1; X[2] = 1; X[1] = 1; X[0] = 1;
			Y[3] = 1; Y[2] = 1; Y[1] = 1; Y[0] = 0;
			Z = 0;
			#10
			
			X[3] = 0; X[2] = 0; X[1] = 1; X[0] = 0;
			Y[3] = 1; Y[2] = 0; Y[1] = 1; Y[0] = 0;
			Z = 1;
			#10
			
			X[3] = 1; X[2] = 1; X[1] = 1; X[0] = 1;
			Y[3] = 0; Y[2] = 1; Y[1] = 1; Y[0] = 1;
			Z = 0;
			#10
			
			X[3] = 0; X[2] = 1; X[1] = 1; X[0] = 0;
			Y[3] = 1; Y[2] = 0; Y[1] = 1; Y[0] = 0;
			Z = 1;
			#10
			
			X[3] = 1; X[2] = 1; X[1] = 0; X[0] = 1;
			Y[3] = 1; Y[2] = 1; Y[1] = 0; Y[0] = 1;
			Z = 1;
			#10
			
			X[3] = 1; X[2] = 0; X[1] = 0; X[0] = 0;
			Y[3] = 0; Y[2] = 1; Y[1] = 1; Y[0] = 0;
			Z = 1;
			#10
			
			X[3] = 1; X[2] = 0; X[1] = 1; X[0] = 0;
			Y[3] = 1; Y[2] = 1; Y[1] = 1; Y[0] = 1;
			Z = 0;
			#10
			
		$finish;
	end
endmodule