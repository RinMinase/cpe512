module tb_fourBitAdder;
	reg [3:0] A, B;
	reg	Cin;
	
	wire [3:0] S;
	wire Cout;
	
	fourBitAdder UUT(A, B, Cin, S, Cout);
	
	initial
		begin
			$dumpfile("fourBitAdder.vpd");
			$dumpvars;

			A[3] = 1; A[2] = 0; A[1] = 1; A[0] = 0;
			B[3] = 0; B[2] = 1; B[1] = 0; B[0] = 1;
			Cin = 0;
			#10
			
			A[3] = 1; A[2] = 1; A[1] = 0; A[0] = 1;
			B[3] = 1; B[2] = 0; B[1] = 0; B[0] = 0;
			Cin = 1;
			#10
			
			A[3] = 0; A[2] = 1; A[1] = 0; A[0] = 0;
			B[3] = 1; B[2] = 1; B[1] = 0; B[0] = 0;
			Cin = 0;
			#10
			
			A[3] = 1; A[2] = 1; A[1] = 1; A[0] = 1;
			B[3] = 1; B[2] = 1; B[1] = 1; B[0] = 0;
			Cin = 0;
			#10
			
			A[3] = 0; A[2] = 0; A[1] = 1; A[0] = 0;
			B[3] = 1; B[2] = 0; B[1] = 1; B[0] = 0;
			Cin = 1;
			#10
			
			A[3] = 1; A[2] = 1; A[1] = 1; A[0] = 1;
			B[3] = 0; B[2] = 1; B[1] = 1; B[0] = 1;
			Cin = 0;
			#10
			
			A[3] = 0; A[2] = 1; A[1] = 1; A[0] = 0;
			B[3] = 1; B[2] = 0; B[1] = 1; B[0] = 0;
			Cin = 1;
			#10
			
			A[3] = 1; A[2] = 1; A[1] = 0; A[0] = 1;
			B[3] = 1; B[2] = 1; B[1] = 0; B[0] = 1;
			Cin = 1;
			#10
			
			A[3] = 1; A[2] = 0; A[1] = 0; A[0] = 0;
			B[3] = 0; B[2] = 1; B[1] = 1; B[0] = 0;
			Cin = 1;
			#10
			
			A[3] = 1; A[2] = 0; A[1] = 1; A[0] = 0;
			B[3] = 1; B[2] = 1; B[1] = 1; B[0] = 1;
			Cin = 0;
			#10
			
		$finish;
	end
endmodule