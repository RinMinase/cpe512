module tb_accumulator;
	reg [3:0] a,b, m;
	reg cin;

	wire [3:0] r;
	wire ovf;

	reg Clk, nReset;

	wire CBF;
	wire [3:0] Y;

	fourBitAluWithShifter UUT (.A(a), .B(b), .Cin(cin), .Mode(m), .R(r), .overFlow(ovf));
	accumulator UUT2({ovf,r},Clk,nReset,CBF,Y);

	initial begin

		$dumpfile("accumulator.vpd");
		$dumpvars;
	end

	initial
		Clk = 0;

	always
		#5 Clk = ~Clk;

	initial begin
		nReset <= 0;
		#10
		nReset <= 1;
	end

	initial begin


a = 4'b1111; b = 4'b1110; cin = 4'b0110; m = 4'b0000; #10 
a = 4'b0100; b = 4'b1110; cin = 4'b1110; m = 4'b0000; #10 
a = 4'b1100; b = 4'b0101; cin = 4'b1111; m = 4'b0000; #10

a = 4'b1001; b = 4'b1101; cin = 4'd1; m = 4'b0001; #10 
a = 4'b0101; b = 4'b1010; cin = 4'd1; m = 4'b0001; #10 
a = 4'b0110; b = 4'b1110; cin = 4'd1; m = 4'b0001; #10 

a = 4'b1110; b = 4'b1011; cin = 4'b0110; m = 4'b0010; #10 
a = 4'b1111; b = 4'b1011; cin = 4'b1010; m = 4'b0010; #10 
a = 4'b1010; b = 4'b0100; cin = 4'b0101; m = 4'b0010; #10 

a = 4'b1010; b = 4'b0101; cin = 4'b0001; m = 4'b0011; #10
a = 4'b1111; b = 4'b1110; cin = 4'b0110; m = 4'b0011; #10 
a = 4'b0100; b = 4'b1110; cin = 4'b1110; m = 4'b0011; #10 

a = 4'b1100; b = 4'b0101; cin = 4'b1111; m = 4'b0100; #10 
a = 4'b1001; b = 4'b1101; cin = 4'b1011; m = 4'b0100; #10 
a = 4'b0101; b = 4'b1010; cin = 4'b0111; m = 4'b0100; #10 

a = 4'b0110; b = 4'b1110; cin = 4'b1001; m = 4'b0101; #10 
a = 4'b1110; b = 4'b1011; cin = 4'b0110; m = 4'b0101; #10 
a = 4'b1111; b = 4'b1011; cin = 4'b1010; m = 4'b0101; #10 

a = 4'b1010; b = 4'b0100; cin = 4'b0101; m = 4'b0110; #10 
a = 4'b1010; b = 4'b0101; cin = 4'b0001; m = 4'b0110; #10
a = 4'b1110; b = 4'b1011; cin = 4'b0110; m = 4'b0110; #10 

a = 4'b1111; b = 4'b1011; cin = 4'b1010; m = 4'b0111; #10 
a = 4'b1010; b = 4'b0100; cin = 4'b0101; m = 4'b0111; #10 
a = 4'b1010; b = 4'b0101; cin = 4'b0001; m = 4'b0111; #10

a = 4'b1111; b = 4'b1110; cin = 4'b0110; m = 4'b1000; #10 
a = 4'b0100; b = 4'b1110; cin = 4'b1110; m = 4'b1000; #10 
a = 4'b1100; b = 4'b0101; cin = 4'b1111; m = 4'b1000; #10

a = 4'b1001; b = 4'b1101; cin = 4'b0110; m = 4'b1001; #10 
a = 4'b0101; b = 4'b1010; cin = 4'b1110; m = 4'b1001; #10 
a = 4'b0110; b = 4'b1110; cin = 4'b1111; m = 4'b1001; #10 

a = 4'b1110; b = 4'b1011; cin = 4'b0110; m = 4'b1010; #10 
a = 4'b1111; b = 4'b1011; cin = 4'b1010; m = 4'b1010; #10 
a = 4'b1010; b = 4'b0100; cin = 4'b0101; m = 4'b1010; #10 

a = 4'b1010; b = 4'b0101; cin = 4'b0001; m = 4'b1011; #10
a = 4'b1111; b = 4'b1110; cin = 4'b0110; m = 4'b1011; #10 
a = 4'b0100; b = 4'b1110; cin = 4'b1110; m = 4'b1011; #10 

a = 4'b1100; b = 4'b0101; cin = 4'b1111; m = 4'b1100; #10 
a = 4'b1001; b = 4'b1101; cin = 4'b1011; m = 4'b1100; #10 
a = 4'b0101; b = 4'b1010; cin = 4'b0111; m = 4'b1100; #10 

a = 4'b0110; b = 4'b1110; cin = 4'b1001; m = 4'b1101; #10 
a = 4'b1110; b = 4'b1011; cin = 4'b0110; m = 4'b1101; #10 
a = 4'b1111; b = 4'b1011; cin = 4'b1010; m = 4'b1101; #10 

a = 4'b1010; b = 4'b0100; cin = 4'b0101; m = 4'b1110; #10 
a = 4'b1010; b = 4'b0101; cin = 4'b0001; m = 4'b1110; #10
a = 4'b1110; b = 4'b1011; cin = 4'b0110; m = 4'b1110; #10 

a = 4'b1111; b = 4'b1011; cin = 4'b1010; m = 4'b1111; #10 
a = 4'b1010; b = 4'b0100; cin = 4'b0101; m = 4'b1111; #10 
a = 4'b1010; b = 4'b0101; cin = 4'b0001; m = 4'b1111; #10



		$finish;

	end

endmodule