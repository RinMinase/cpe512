module tb_fourBitSubtractor;
	reg [3:0] A, B;
	
	wire [3:0] D;
	wire Bout;
	
	fourBitSubtractor UUT(A, B, D, Bout);
	
	initial
		begin
			$dumpfile("fourBitSubtractor.vpd");
			$dumpvars;
			
			A[3] = 1; A[2] = 0; A[1] = 1; A[0] = 0;
			B[3] = 0; B[2] = 1; B[1] = 0; B[0] = 1;
			#10
			
			A[3] = 1; A[2] = 1; A[1] = 0; A[0] = 1;
			B[3] = 1; B[2] = 0; B[1] = 0; B[0] = 0;
			#10
			
			A[3] = 0; A[2] = 1; A[1] = 0; A[0] = 0;
			B[3] = 1; B[2] = 1; B[1] = 0; B[0] = 0;
			#10
			
			A[3] = 1; A[2] = 1; A[1] = 1; A[0] = 1;
			B[3] = 1; B[2] = 1; B[1] = 1; B[0] = 0;
			#10
			
			A[3] = 0; A[2] = 0; A[1] = 1; A[0] = 0;
			B[3] = 1; B[2] = 0; B[1] = 1; B[0] = 0;
			#10
			
			A[3] = 1; A[2] = 1; A[1] = 1; A[0] = 1;
			B[3] = 0; B[2] = 1; B[1] = 1; B[0] = 1;
			#10
			
			A[3] = 0; A[2] = 1; A[1] = 1; A[0] = 0;
			B[3] = 1; B[2] = 0; B[1] = 1; B[0] = 0;
			#10
			
			A[3] = 1; A[2] = 1; A[1] = 0; A[0] = 1;
			B[3] = 1; B[2] = 1; B[1] = 0; B[0] = 1;
			#10
			
			A[3] = 1; A[2] = 0; A[1] = 0; A[0] = 0;
			B[3] = 0; B[2] = 1; B[1] = 1; B[0] = 0;
			#10
			
			A[3] = 1; A[2] = 0; A[1] = 1; A[0] = 0;
			B[3] = 1; B[2] = 1; B[1] = 1; B[0] = 1;
			#10
			
		$finish;
	end
endmodule